module hello;
initial begin;
    $display("hello learncocotb.com");
end
endmodule
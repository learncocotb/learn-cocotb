module hello;
initial begin;
    $display("hello learncocotb.com ayyyyyy");
end
endmodule